//-- Verilog hello world example
//-  A NOT gate
module inv(input A, output B);
wire A;
wire B;


  assign B = !A;

endmodule


